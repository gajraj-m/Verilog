`include "CLA_16bit.v"

module q2_tb;
    reg [15:0] A,B;
    reg C_In;
    wire [15:0] Sum;
    wire c_out;

    CLA_16bit inst0(c_out, Sum, A, B, C_In);

    initial begin

        $monitor("%t| A = %d, B = %d, C_In = %b | C_Out = %b | Sum = %d", $time, A, B, C_In, c_out, Sum);

        A = 16'b0000000000010000; B = 16'b0000000010000000; C_In = 1'b1;
        #1 A = 16'b0000001000000000; B = 16'b0000010000110001; C_In = 1'b1;
        #1 A = 16'b1000000001000000; B = 16'b0000000000000101; C_In = 1'b0;
        #1 A = 16'b0000000001100100; B = 16'b0000000000001000; C_In = 1'b0;
        #1 A = 16'b0000010011000000; B = 16'b0000000011100001; C_In = 1'b1;
        #1 A = 16'b1000010000000000; B = 16'b0001100000000000; C_In = 1'b0;
        #1 A = 16'b0010110000000000; B = 16'b0010000010010100; C_In = 1'b1;
        #1 A = 16'b1000000000000110; B = 16'b1100010000100001; C_In = 1'b0;
    end

endmodule