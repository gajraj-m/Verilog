module xor_gate(output c, input a, b);

xor(c, a, b);

endmodule